module first (
	input wire switch,
	output wire led
);
assign led = switch;

endmodule
